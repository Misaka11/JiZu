module mips(clk,rst);
	input clk;
	input rst;
	datapath _dp(clk,rst);
endmodule